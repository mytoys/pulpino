
module boot_code
(
    input  logic        CLK,
    input  logic        RSTN,

    input  logic        CSN,
    input  logic [9:0]  A,
    output logic [31:0] Q
  );

  const logic [0:547] [31:0] mem = {
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h0100006F,
    32'h0100006F,
    32'h0080006F,
    32'h0040006F,
    32'h0000006F,
    32'h00000093,
    32'h00008113,
    32'h00008193,
    32'h00008213,
    32'h00008293,
    32'h00008313,
    32'h00008393,
    32'h00008413,
    32'h00008493,
    32'h00008513,
    32'h00008593,
    32'h00008613,
    32'h00008693,
    32'h00008713,
    32'h00008793,
    32'h00008813,
    32'h00008893,
    32'h00008913,
    32'h00008993,
    32'h00008A13,
    32'h00008A93,
    32'h00008B13,
    32'h00008B93,
    32'h00008C13,
    32'h00008C93,
    32'h00008D13,
    32'h00008D93,
    32'h00008E13,
    32'h00008E93,
    32'h00008F13,
    32'h00008F93,
    32'h00100117,
    32'hEF410113,
    32'h00000D17,
    32'h748D0D13,
    32'h00000D97,
    32'h744D8D93,
    32'h01BD5863,
    32'h000D2023,
    32'h004D0D13,
    32'hFFADDCE3,
    32'h00000513,
    32'h00000593,
    32'h014000EF,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h4505715D,
    32'hC4A2C686,
    32'hC0CAC2A6,
    32'hDC52DE4E,
    32'hD85ADA56,
    32'hD462D65E,
    32'hD06AD266,
    32'h244000EF,
    32'h45014585,
    32'h448000EF,
    32'h87936785,
    32'h0001BB87,
    32'hFFF517FD,
    32'h27B74711,
    32'h85371A10,
    32'hC3D80000,
    32'h051345C5,
    32'h00EF6A45,
    32'h46814760,
    32'h45A14601,
    32'h00EF4519,
    32'h45012C20,
    32'h310000EF,
    32'h458164C1,
    32'h00EF4505,
    32'h14FD33E0,
    32'h00EF4405,
    32'h8D653660,
    32'hFE851DE3,
    32'h85B646A1,
    32'h05F00613,
    32'h06100513,
    32'h294000EF,
    32'h00EF4501,
    32'h64C12E20,
    32'h85224581,
    32'h310000EF,
    32'h00EF14FD,
    32'h8D6533A0,
    32'hFE851DE3,
    32'h45214581,
    32'h2A8000EF,
    32'h02000693,
    32'h40000637,
    32'h051345A1,
    32'h00EF0EB0,
    32'h051325E0,
    32'h00EF1000,
    32'h45812AA0,
    32'h00EF4509,
    32'h05932DA0,
    32'h850A1000,
    32'h31C000EF,
    32'h00008537,
    32'h45D54CB2,
    32'h6B850513,
    32'h4C124982,
    32'h4BD24942,
    32'h00EF4B72,
    32'h45813D20,
    32'h00EF4521,
    32'h5E6325A0,
    32'h64A10790,
    32'h0C334401,
    32'h8AB7413C,
    32'h84930000,
    32'h8A377144,
    32'h6D050000,
    32'h00899613,
    32'h02000693,
    32'h051345A1,
    32'h00EF0EB0,
    32'h65211F60,
    32'h244000EF,
    32'h45094581,
    32'h274000EF,
    32'h013C0533,
    32'h00EF65A1,
    32'h45992B60,
    32'h6D0A8513,
    32'h37C000EF,
    32'h00445513,
    32'h95264585,
    32'h370000EF,
    32'h00F47513,
    32'h95264585,
    32'h364000EF,
    32'h45990405,
    32'h6D8A0513,
    32'h358000EF,
    32'h00EF99EA,
    32'h91E338E0,
    32'h6441FA8C,
    32'h4485147D,
    32'h258000EF,
    32'h1DE38D61,
    32'h8537FE95,
    32'h45B50000,
    32'h6E050513,
    32'h330000EF,
    32'h368000EF,
    32'h45214581,
    32'h1B4000EF,
    32'h07605E63,
    32'h440164A1,
    32'h00008AB7,
    32'h71448493,
    32'h00008A37,
    32'h412B8BB3,
    32'h16136985,
    32'h06930089,
    32'h45A10200,
    32'h0EB00513,
    32'h150000EF,
    32'h00EF6521,
    32'h458119E0,
    32'h00EF4509,
    32'h85331CE0,
    32'h65A1012B,
    32'h210000EF,
    32'h85134599,
    32'h00EF6D0A,
    32'h55132D60,
    32'h45850044,
    32'h00EF9526,
    32'h75132CA0,
    32'h458500F4,
    32'h00EF9526,
    32'h04052BE0,
    32'h05134599,
    32'h00EF6D8A,
    32'h994E2B20,
    32'h2E8000EF,
    32'hFA8B11E3,
    32'h00008537,
    32'h6F050513,
    32'h02200593,
    32'h298000EF,
    32'h2D0000EF,
    32'h1A107737,
    32'h00072423,
    32'h08000793,
    32'h2E236725,
    32'h978284F7,
    32'h450140B6,
    32'h44964426,
    32'h59F24906,
    32'h5AD25A62,
    32'h5BB25B42,
    32'h5C925C22,
    32'h61615D02,
    32'h00008082,
    32'hFF010113,
    32'h00812423,
    32'h00000593,
    32'h00050413,
    32'h00F00513,
    32'h00112623,
    32'h00912223,
    32'h290000EF,
    32'h00000593,
    32'h00E00513,
    32'h284000EF,
    32'h00000593,
    32'h00D00513,
    32'h278000EF,
    32'h00000593,
    32'h00C00513,
    32'h26C000EF,
    32'h04805E63,
    32'h00100493,
    32'h00000593,
    32'h01000513,
    32'h258000EF,
    32'h04940463,
    32'h00000593,
    32'h00B00513,
    32'h248000EF,
    32'h00200793,
    32'h02F40A63,
    32'h00000593,
    32'h00000513,
    32'h234000EF,
    32'h00300793,
    32'h02F40063,
    32'h00048513,
    32'h00C12083,
    32'h00812403,
    32'h00412483,
    32'h00000593,
    32'h01010113,
    32'h2100006F,
    32'h00C12083,
    32'h00812403,
    32'h00412483,
    32'h01010113,
    32'h00008067,
    32'h00004737,
    32'hF0070713,
    32'h00869693,
    32'h02000793,
    32'h40B787B3,
    32'h00E6F6B3,
    32'h03F5F593,
    32'h1A102737,
    32'h00F51533,
    32'h00B6E5B3,
    32'h00A72423,
    32'h00C72623,
    32'h00B72823,
    32'h00008067,
    32'h01051513,
    32'h01059593,
    32'h01055513,
    32'h00A5E5B3,
    32'h1A1027B7,
    32'h00B7AA23,
    32'h00008067,
    32'h1A102737,
    32'h01072783,
    32'hFF010113,
    32'h00F12623,
    32'h00C12783,
    32'h01051513,
    32'h01079793,
    32'h0107D793,
    32'h00F56533,
    32'h00A12623,
    32'h00C12783,
    32'h01010113,
    32'h00F72823,
    32'h00008067,
    32'h00100793,
    32'h00858593,
    32'h00B795B3,
    32'h00A79533,
    32'h000017B7,
    32'hF0078793,
    32'h00F5F5B3,
    32'h0FF57513,
    32'h00A5E533,
    32'h1A1027B7,
    32'h00A7A023,
    32'h00008067,
    32'h1A1027B7,
    32'h0007A783,
    32'hFF010113,
    32'h00F12623,
    32'h00C12503,
    32'h01010113,
    32'h00008067,
    32'h4055D793,
    32'hFF010113,
    32'h7FF7F793,
    32'h01F5F593,
    32'h00F12423,
    32'h00058863,
    32'h00812783,
    32'h00178793,
    32'h00F12423,
    32'h00012623,
    32'h00C12683,
    32'h00812783,
    32'h1A102737,
    32'h00070813,
    32'h04F6D063,
    32'h00072783,
    32'h4107D793,
    32'h0FF7F793,
    32'hFE078AE3,
    32'h00C12783,
    32'h02082583,
    32'h00C12683,
    32'h00279793,
    32'h00168693,
    32'h00D12623,
    32'h00C12603,
    32'h00812683,
    32'h00F507B3,
    32'h00B7A023,
    32'hFCD644E3,
    32'h01010113,
    32'h00008067,
    32'h1A1076B7,
    32'h0046A703,
    32'h1A1007B7,
    32'h00276713,
    32'h00E6A223,
    32'h08300713,
    32'h00E7A623,
    32'h0085D613,
    32'h0A700713,
    32'h0FF5F593,
    32'h00C7A223,
    32'h00B7A023,
    32'h00E7A423,
    32'h00300713,
    32'h00E7A623,
    32'h0047A703,
    32'h0F077713,
    32'h00276713,
    32'h00E7A223,
    32'h00008067,
    32'h1A100737,
    32'h02058A63,
    32'h04050613,
    32'h01472783,
    32'h0207F793,
    32'hFE078CE3,
    32'h00150513,
    32'hFFF54683,
    32'h1A1007B7,
    32'hFFF58593,
    32'h00D7A023,
    32'hFCC50CE3,
    32'hFC059EE3,
    32'h00008067,
    32'h00008067,
    32'h1A100737,
    32'h01472783,
    32'h0407F793,
    32'hFE078CE3,
    32'h00008067,
    32'h1A1076B7,
    32'h0006A783,
    32'hFF010113,
    32'h00F12623,
    32'h00100793,
    32'h00C12703,
    32'h00A797B3,
    32'hFFF7C793,
    32'h00E7F7B3,
    32'h00F12623,
    32'h00C12783,
    32'h00A595B3,
    32'h00F5E533,
    32'h00A12623,
    32'h00C12783,
    32'h01010113,
    32'h00F6A023,
    32'h00008067,
    32'h64616F4C,
    32'h20676E69,
    32'h6D6F7266,
    32'h49505320,
    32'h0000000A,
    32'h79706F43,
    32'h20676E69,
    32'h74736E49,
    32'h74637572,
    32'h736E6F69,
    32'h0000000A,
    32'h636F6C42,
    32'h0000206B,
    32'h6E6F6420,
    32'h00000A65,
    32'h79706F43,
    32'h20676E69,
    32'h61746144,
    32'h0000000A,
    32'h656E6F44,
    32'h756A202C,
    32'h6E69706D,
    32'h6F742067,
    32'h736E4920,
    32'h63757274,
    32'h6E6F6974,
    32'h4D415220,
    32'h00000A2E,
    32'h33323130,
    32'h37363534,
    32'h42413938,
    32'h46454443,
    32'h00000010,
    32'h00000000,
    32'h00527A01,
    32'h01010401,
    32'h00020D1B,
    32'h00000038,
    32'h00000018,
    32'hFFFFFA10,
    32'h0000025E,
    32'h500E4200,
    32'h7F01115A,
    32'h117E0811,
    32'h12117D09,
    32'h7B13117C,
    32'h117A1411,
    32'h16117915,
    32'h77171178,
    32'h11761811,
    32'h1A117519,
    32'h00000074,
    32'h0000001C,
    32'h00000054,
    32'hFFFFFC34,
    32'h000000B4,
    32'h100E4400,
    32'h7E081148,
    32'h7F011150,
    32'h007D0911,
    32'h00000010,
    32'h00000074,
    32'hFFFFFCC8,
    32'h00000038,
    32'h00000000,
    32'h00000010,
    32'h00000088,
    32'hFFFFFCEC,
    32'h0000001C,
    32'h00000000,
    32'h00000010,
    32'h0000009C,
    32'hFFFFFCF4,
    32'h00000038,
    32'h100E4C00,
    32'h00000010,
    32'h000000B0,
    32'hFFFFFD18,
    32'h00000030,
    32'h00000000,
    32'h00000010,
    32'h000000C4,
    32'hFFFFFD34,
    32'h0000001C,
    32'h100E4C00,
    32'h00000010,
    32'h000000D8,
    32'hFFFFFD3C,
    32'h00000080,
    32'h100E4800,
    32'h00000010,
    32'h000000EC,
    32'hFFFFFDA8,
    32'h00000050,
    32'h00000000,
    32'h00000010,
    32'h00000100,
    32'hFFFFFDE4,
    32'h0000003C,
    32'h00000000,
    32'h00000010,
    32'h00000114,
    32'hFFFFFE0C,
    32'h00000014,
    32'h00000000,
    32'h00000010,
    32'h00000128,
    32'hFFFFFE0C,
    32'h00000048,
    32'h100E4C00,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000};

  logic [9:0] A_Q;

  always_ff @(posedge CLK, negedge RSTN)
  begin
    if (~RSTN)
      A_Q <= '0;
    else
      if (~CSN)
        A_Q <= A;
  end

  assign Q = mem[A_Q];

endmodule